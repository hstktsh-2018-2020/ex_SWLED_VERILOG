`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:55:37 12/12/2017 
// Design Name: 
// Module Name:    ex_SWLED_VERILOG 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ex_SWLED_VERILOG(
    input CLK,
    output LED0
    );

assign LED0 = CLK;

endmodule

